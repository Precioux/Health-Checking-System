/*--  *******************************************************
--  Computer Architecture Course, Laboratory Sources 
--  Amirkabir University of Technology (Tehran Polytechnic)
--  Department of Computer Engineering (CE-AUT)
--  https://ce[dot]aut[dot]ac[dot]ir
--  *******************************************************
--  All Rights reserved (C) 2020-2021
--  *******************************************************
--  Student ID  : 9833016              9839039
--  Student Name: Amirhossein Poolad & Samin Mahdipour
--  Student Mail: 
--  *******************************************************
--  Additional Comments:
--
--*/

/*-----------------------------------------------------------
---  Module Name: Temperature Analyzer
-----------------------------------------------------------*/
`timescale 1ns / 1ps
module tb_temperatureAnalyzer();
reg [7:0] t;
wire ht;
wire lt;
temperatureAnalyzer a(t,ht,lt);
initial 
    begin 
	  t=7'b0000000;
	  #10;
	  t=7'b0000001;
	  #10;
	  t=7'b0000010;
	  #10;
	  t=7'b0000011;
	  #10;
	  t=7'b0000100;
	  #10;
	  t=7'b0000101;
	  #10;
	  t=7'b0000110;
	  #10;
	  t=7'b0000111;
	  #10;
	  t=7'b0001000;
	  #10;
	  t=7'b0001001;
	  #10;
	  t=7'b0001010;
	  #10;
	  t=7'b0001011;
	  #10;
	  t=7'b0001100;
	  #10;
	  t=7'b0001101;
	  #10;
	  t=7'b0001110;
	  #10;
	  t=7'b0001111;
	  #10;
     t=7'b0010000;
	  #10;
	  t=7'b0010001;
	  #10;
	  t=7'b0010010;
	  #10;
	  t=7'b0010011;
	  #10;
	  t=7'b0010100;
	  #10;
	  t=7'b0010101;
	  #10;
	  t=7'b0010110;
	  #10;
	  t=7'b0010111;
	  #10;
	  t=7'b0011000;
	  #10;
	  t=7'b0011001;
	  #10;
	  t=7'b0011010;
	  #10;
	  t=7'b0011011;
	  #10;
	  t=7'b0011100;
	  #10;
	  t=7'b0011101;
	  #10;
	  t=7'b0011110;
	  #10;
	  t=7'b0011111;
	  #10;
	  t=7'b0100000;
	  #10;
	  t=7'b0100001;
	  #10;
	  t=7'b0100010;
	  #10;
	  t=7'b0100011;
	  #10;
	  t=7'b0100100;
	  #10;
	  t=7'b0100101;
	  #10;
	  t=7'b0100110;
	  #10;
	  t=7'b0100111;
	  #10;
	  t=7'b0101000;
	  #10;
	  t=7'b0101001;
	  #10;
	  t=7'b0101010;
	  #10;
	  t=7'b0101011;
	  #10;
	  t=7'b0101100;
	  #10;
	  t=7'b0101101;
	  #10;
	  t=7'b0101110;
	  #10;
	  t=7'b0101111;
	  #10;
     t=7'b0110000;
	  #10;
	  t=7'b0110001;
	  #10;
	  t=7'b0110010;
	  #10;
	  t=7'b0110011;
	  #10;
	  t=7'b0110100;
	  #10;
	  t=7'b0110101;
	  #10;
	  t=7'b0110110;
	  #10;
	  t=7'b0110111;
	  #10;
	  t=7'b0111000;
	  #10;
	  t=7'b0111001;
	  #10;
	  t=7'b0111010;
	  #10;
	  t=7'b0111011;
	  #10;
	  t=7'b0111100;
	  #10;
	  t=7'b0111101;
	  #10;
	  t=7'b0111110;
	  #10;
	  t=7'b0111111;
	  #10;
	  t=7'b1000000;
	  #10;
	  t=7'b1000001;
	  #10;
	  t=7'b1000010;
	  #10;
	  t=7'b1000011;
	  #10;
	  t=7'b1000100;
	  #10;
	  t=7'b1000101;
	  #10;
	  t=7'b1000110;
	  #10;
	  t=7'b1000111;
	  #10;
	  t=7'b1001000;
	  #10;
	  t=7'b1001001;
	  #10;
	  t=7'b1001010;
	  #10;
	  t=7'b1001011;
	  #10;
	  t=7'b1001100;
	  #10;
	  t=7'b1001101;
	  #10;
	  t=7'b1001110;
	  #10;
	  t=7'b1001111;
	  #10;
     t=7'b1010000;
	  #10;
	  t=7'b1010001;
	  #10;
	  t=7'b1010010;
	  #10;
	  t=7'b1010011;
	  #10;
	  t=7'b1010100;
	  #10;
	  t=7'b1010101;
	  #10;
	  t=7'b1010110;
	  #10;
	  t=7'b1010111;
	  #10;
	  t=7'b1011000;
	  #10;
	  t=7'b1011001;
	  #10;
	  t=7'b1011010;
	  #10;
	  t=7'b1011011;
	  #10;
	  t=7'b1011100;
	  #10;
	  t=7'b1011101;
	  #10;
	  t=7'b1011110;
	  #10;
	  t=7'b1011111;
	  #10;
	  t=7'b1100000;
	  #10;
	  t=7'b1100001;
	  #10;
	  t=7'b1100010;
	  #10;
	  t=7'b1100011;
	  #10;
	  t=7'b1100100;
	  #10;
	  t=7'b1100101;
	  #10;
	  t=7'b1100110;
	  #10;
	  t=7'b1100111;
	  #10;
	  t=7'b1101000;
	  #10;
	  t=7'b1101001;
	  #10;
	  t=7'b1101010;
	  #10;
	  t=7'b1101011;
	  #10;
	  t=7'b1101100;
	  #10;
	  t=7'b1101101;
	  #10;
	  t=7'b1101110;
	  #10;
	  t=7'b1101111;
	  #10;
     t=7'b1110000;
	  #10;
	  t=7'b1110001;
	  #10;
	  t=7'b1110010;
	  #10;
	  t=7'b1110011;
	  #10;
	  t=7'b1110100;
	  #10;
	  t=7'b1110101;
	  #10;
	  t=7'b1110110;
	  #10;
	  t=7'b1110111;
	  #10;
	  t=7'b1111000;
	  #10;
	  t=7'b1111001;
	  #10;
	  t=7'b1111010;
	  #10;
	  t=7'b1111011;
	  #10;
	  t=7'b1111100;
	  #10;
	  t=7'b1111101;
	  #10;
	  t=7'b1111110;
	  #10;
	  t=7'b1111111;
	 end
	endmodule
module temperatureAnalyzer(
 temperature,
 highTempAbnormality,
  lowTempAbnormality
 );
input [7:0] temperature;
output lowTempAbnormality;
output highTempAbnormality;
 assign lowTempAbnormality = (temperature < 35);
 assign highTempAbnormality = (temperature > 39);
endmodule
