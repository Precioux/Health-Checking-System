/*--  *******************************************************
--  Computer Architecture Course, Laboratory Sources 
--  Amirkabir University of Technology (Tehran Polytechnic)
--  Department of Computer Engineering (CE-AUT)
--  https://ce[dot]aut[dot]ac[dot]ir
--  *******************************************************
--  All Rights reserved (C) 2020-2021
--  *******************************************************
--  Student ID  : 9833016              9839039
--  Student Name: Amirhossein Poolad & Samin Mahdipour
--  Student Mail: 
--  *******************************************************
--  Additional Comments:
--
--*/

/*-----------------------------------------------------------
---  Module Name: 4 Bit Ripple Carry Adder
-----------------------------------------------------------*/
`timescale 1ns / 1ps
module tb_ripple_carry_adder();
reg [3:0]a;
reg [3:0]b;
wire c;
wire [3:0]s;
initial 
    begin 
        a=4'b0000;
        #10;
        b=4'b0000;
        #10;
        b=4'b0001;
        #10;
        b=4'b0010;
        #10;
        b=4'b0011;
        #10;
        b=4'b0100;
        #10;
        b=4'b0101;
        #10;
        b=4'b0110;
        #10;
        b=4'b0111;
        #10;
        b=4'b1000;
        #10;
        b=4'b1001;
        #10;
        b=4'b1010;
        #10;
        b=4'b1011;
        #10;
        b=4'b1100;
        #10;
        b=4'b1101;
        #10;
        b=4'b1110;
        #10;
        b=4'b1111;
        #10;
        a=4'b0001;
         #10;
        b=4'b0000;
        #10;
        b=4'b0001;
        #10;
        b=4'b0010;
        #10;
        b=4'b0011;
        #10;
        b=4'b0100;
        #10;
        b=4'b0101;
        #10;
        b=4'b0110;
        #10;
        b=4'b0111;
        #10;
        b=4'b1000;
        #10;
        b=4'b1001;
        #10;
        b=4'b1010;
        #10;
        b=4'b1011;
        #10;
        b=4'b1100;
        #10;
        b=4'b1101;
        #10;
        b=4'b1110;
        #10;
        b=4'b1111;
        #10;
        a=4'b0010;
         #10;
        b=4'b0000;
        #10;
        b=4'b0001;
        #10;
        b=4'b0010;
        #10;
        b=4'b0011;
        #10;
        b=4'b0100;
        #10;
        b=4'b0101;
        #10;
        b=4'b0110;
        #10;
        b=4'b0111;
        #10;
        b=4'b1000;
        #10;
        b=4'b1001;
        #10;
        b=4'b1010;
        #10;
        b=4'b1011;
        #10;
        b=4'b1100;
        #10;
        b=4'b1101;
        #10;
        b=4'b1110;
        #10;
        b=4'b1111;
        #10;
        a=4'b0011;
         #10;
        b=4'b0000;
        #10;
        b=4'b0001;
        #10;
        b=4'b0010;
        #10;
        b=4'b0011;
        #10;
        b=4'b0100;
        #10;
        b=4'b0101;
        #10;
        b=4'b0110;
        #10;
        b=4'b0111;
        #10;
        b=4'b1000;
        #10;
        b=4'b1001;
        #10;
        b=4'b1010;
        #10;
        b=4'b1011;
        #10;
        b=4'b1100;
        #10;
        b=4'b1101;
        #10;
        b=4'b1110;
        #10;
        b=4'b1111;
        #10;
        a=4'b0100;
         #10;
        b=4'b0000;
        #10;
        b=4'b0001;
        #10;
        b=4'b0010;
        #10;
        b=4'b0011;
        #10;
        b=4'b0100;
        #10;
        b=4'b0101;
        #10;
        b=4'b0110;
        #10;
        b=4'b0111;
        #10;
        b=4'b1000;
        #10;
        b=4'b1001;
        #10;
        b=4'b1010;
        #10;
        b=4'b1011;
        #10;
        b=4'b1100;
        #10;
        b=4'b1101;
        #10;
        b=4'b1110;
        #10;
        b=4'b1111;
        #10;
        a=4'b0101;
         #10;
        b=4'b0000;
        #10;
        b=4'b0001;
        #10;
        b=4'b0010;
        #10;
        b=4'b0011;
        #10;
        b=4'b0100;
        #10;
        b=4'b0101;
        #10;
        b=4'b0110;
        #10;
        b=4'b0111;
        #10;
        b=4'b1000;
        #10;
        b=4'b1001;
        #10;
        b=4'b1010;
        #10;
        b=4'b1011;
        #10;
        b=4'b1100;
        #10;
        b=4'b1101;
        #10;
        b=4'b1110;
        #10;
        b=4'b1111;
        #10;
        a=4'b0110;
         #10;
        b=4'b0000;
        #10;
        b=4'b0001;
        #10;
        b=4'b0010;
        #10;
        b=4'b0011;
        #10;
        b=4'b0100;
        #10;
        b=4'b0101;
        #10;
        b=4'b0110;
        #10;
        b=4'b0111;
        #10;
        b=4'b1000;
        #10;
        b=4'b1001;
        #10;
        b=4'b1010;
        #10;
        b=4'b1011;
        #10;
        b=4'b1100;
        #10;
        b=4'b1101;
        #10;
        b=4'b1110;
        #10;
        b=4'b1111;
        #10;
        a=4'b0111;
         #10;
        b=4'b0000;
        #10;
        b=4'b0001;
        #10;
        b=4'b0010;
        #10;
        b=4'b0011;
        #10;
        b=4'b0100;
        #10;
        b=4'b0101;
        #10;
        b=4'b0110;
        #10;
        b=4'b0111;
        #10;
        b=4'b1000;
        #10;
        b=4'b1001;
        #10;
        b=4'b1010;
        #10;
        b=4'b1011;
        #10;
        b=4'b1100;
        #10;
        b=4'b1101;
        #10;
        b=4'b1110;
        #10;
        b=4'b1111;
        #10;
        a=4'b1000;
         #10;
        b=4'b0000;
        #10;
        b=4'b0001;
        #10;
        b=4'b0010;
        #10;
        b=4'b0011;
        #10;
        b=4'b0100;
        #10;
        b=4'b0101;
        #10;
        b=4'b0110;
        #10;
        b=4'b0111;
        #10;
        b=4'b1000;
        #10;
        b=4'b1001;
        #10;
        b=4'b1010;
        #10;
        b=4'b1011;
        #10;
        b=4'b1100;
        #10;
        b=4'b1101;
        #10;
        b=4'b1110;
        #10;
        b=4'b1111;
        #10;
        a=4'b1001;
         #10;
        b=4'b0000;
        #10;
        b=4'b0001;
        #10;
        b=4'b0010;
        #10;
        b=4'b0011;
        #10;
        b=4'b0100;
        #10;
        b=4'b0101;
        #10;
        b=4'b0110;
        #10;
        b=4'b0111;
        #10;
        b=4'b1000;
        #10;
        b=4'b1001;
        #10;
        b=4'b1010;
        #10;
        b=4'b1011;
        #10;
        b=4'b1100;
        #10;
        b=4'b1101;
        #10;
        b=4'b1110;
        #10;
        b=4'b1111;
        #10;
        a=4'b1010;
         #10;
        b=4'b0000;
        #10;
        b=4'b0001;
        #10;
        b=4'b0010;
        #10;
        b=4'b0011;
        #10;
        b=4'b0100;
        #10;
        b=4'b0101;
        #10;
        b=4'b0110;
        #10;
        b=4'b0111;
        #10;
        b=4'b1000;
        #10;
        b=4'b1001;
        #10;
        b=4'b1010;
        #10;
        b=4'b1011;
        #10;
        b=4'b1100;
        #10;
        b=4'b1101;
        #10;
        b=4'b1110;
        #10;
        b=4'b1111;
        #10;
        a=4'b1011;
         #10;
        b=4'b0000;
        #10;
        b=4'b0001;
        #10;
        b=4'b0010;
        #10;
        b=4'b0011;
        #10;
        b=4'b0100;
        #10;
        b=4'b0101;
        #10;
        b=4'b0110;
        #10;
        b=4'b0111;
        #10;
        b=4'b1000;
        #10;
        b=4'b1001;
        #10;
        b=4'b1010;
        #10;
        b=4'b1011;
        #10;
        b=4'b1100;
        #10;
        b=4'b1101;
        #10;
        b=4'b1110;
        #10;
        b=4'b1111;
        #10;
        a=4'b1100;
         #10;
        b=4'b0000;
        #10;
        b=4'b0001;
        #10;
        b=4'b0010;
        #10;
        b=4'b0011;
        #10;
        b=4'b0100;
        #10;
        b=4'b0101;
        #10;
        b=4'b0110;
        #10;
        b=4'b0111;
        #10;
        b=4'b1000;
        #10;
        b=4'b1001;
        #10;
        b=4'b1010;
        #10;
        b=4'b1011;
        #10;
        b=4'b1100;
        #10;
        b=4'b1101;
        #10;
        b=4'b1110;
        #10;
        b=4'b1111;
        #10;
        a=4'b1101;
         #10;
        b=4'b0000;
        #10;
        b=4'b0001;
        #10;
        b=4'b0010;
        #10;
        b=4'b0011;
        #10;
        b=4'b0100;
        #10;
        b=4'b0101;
        #10;
        b=4'b0110;
        #10;
        b=4'b0111;
        #10;
        b=4'b1000;
        #10;
        b=4'b1001;
        #10;
        b=4'b1010;
        #10;
        b=4'b1011;
        #10;
        b=4'b1100;
        #10;
        b=4'b1101;
        #10;
        b=4'b1110;
        #10;
        b=4'b1111;
        #10;
        a=4'b1110;
         #10;
        b=4'b0000;
        #10;
        b=4'b0001;
        #10;
        b=4'b0010;
        #10;
        b=4'b0011;
        #10;
        b=4'b0100;
        #10;
        b=4'b0101;
        #10;
        b=4'b0110;
        #10;
        b=4'b0111;
        #10;
        b=4'b1000;
        #10;
        b=4'b1001;
        #10;
        b=4'b1010;
        #10;
        b=4'b1011;
        #10;
        b=4'b1100;
        #10;
        b=4'b1101;
        #10;
        b=4'b1110;
        #10;
        b=4'b1111;
        #10;
        a=4'b1111;
         #10;
        b=4'b0000;
        #10;
        b=4'b0001;
        #10;
        b=4'b0010;
        #10;
        b=4'b0011;
        #10;
        b=4'b0100;
        #10;
        b=4'b0101;
        #10;
        b=4'b0110;
        #10;
        b=4'b0111;
        #10;
        b=4'b1000;
        #10;
        b=4'b1001;
        #10;
        b=4'b1010;
        #10;
        b=4'b1011;
        #10;
        b=4'b1100;
        #10;
        b=4'b1101;
        #10;
        b=4'b1110;
        #10;
        b=4'b1111;
        #10;
        $finish;
     end
  endmodule
module ripple_carry_adder(S, C, A, B);
   output [3:0] S; 
   output 	C;  
   input [3:0] 	A;  
   input [3:0] 	B;  

   wire 	C0; 
   wire 	C1;
   wire 	C2; 
	
   full_adder fa0(S[0], C0, A[0], B[0], 0);    
   full_adder fa1(S[1], C1, A[1], B[1], C0);
   full_adder fa2(S[2], C2, A[2], B[2], C1);
   full_adder fa3(S[3], C, A[3], B[3], C2);   
endmodule
