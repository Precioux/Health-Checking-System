`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    01:06:47 07/23/2021 
// Design Name: 
// Module Name:    tb_HealthcareSystemPhase1 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module tb_HealthcareSystemPhase1(
    );

reg [5:0] pressureData;
reg [3:0] bloodPH;
reg [2:0] bloodType;
reg [7:0] fdSensorValue;
reg [7:0] fdFactoryValue;
reg [7:0] bloodSensor;
reg [4:0] factotyBaseTemp;
reg [3:0] factotyTempCoef;
reg [3:0] tempSensorValue;
wire presureAbnormality;
wire bloodAbnormality;
wire fallDetected;
wire [3:0] glycemicIndex;
wire lowTempAbnormality;
wire highTempAbnormality;	 

HealthcareSystemPhase1 hcs(
 pressureData,
 bloodPH,
 bloodType,
 fdSensorValue,
 fdFactoryValue,
 bloodSensor,
 factotyBaseTemp,
 factotyTempCoef,
 tempSensorValue,
 presureAbnormality,
 bloodAbnormality,
 fallDetected,
 glycemicIndex,
 lowTempAbnormality,
 highTempAbnormality);
 
 initial
	begin
	  pressureData=6'b000000;
	  #10;
	  pressureData=6'b000001;
	  #10;
	  pressureData=6'b000010;
	  #10;
	  pressureData=6'b000011;
	  #10;
	  pressureData=6'b000100;
	  #10;
	  pressureData=6'b000101;
	  #10;
	  pressureData=6'b000110;
	  #10;
	  pressureData=6'b000111;
	  #10;
	  pressureData=6'b001000;
	  #10;
	  pressureData=6'b001001;
	  #10;
	  pressureData=6'b001010;
	  #10;
	  pressureData=6'b001011;
	  #10;
	  pressureData=6'b001100;
	  #10;
	  pressureData=6'b001101;
	  #10;
	  pressureData=6'b001110;
	  #10;
	  pressureData=6'b001111;
	  #10;
	  pressureData=6'b010000;
	  #10;
	  pressureData=6'b010001;
	  #10;
	  pressureData=6'b010010;
	  #10;
	  pressureData=6'b010011;
	  #10;
	  pressureData=6'b010100;
	  #10;
	  pressureData=6'b010101;
	  #10;
	  pressureData=6'b010110;
	  #10;
	  pressureData=6'b010111;
	  #10;
	  pressureData=6'b011000;
	  #10;
	  pressureData=6'b011001;
	  #10;
	  pressureData=6'b011010;
	  #10;
	  pressureData=6'b011011;
	  #10;
	  pressureData=6'b011100;
	  #10;
	  pressureData=6'b011101;
	  #10;
	  pressureData=6'b011110;
	  #10;
	  pressureData=6'b011111;
	  #10;
	  pressureData=6'b100000;
	  #10;
	  pressureData=6'b100001;
	  #10;
	  pressureData=6'b100010;
	  #10;
	  pressureData=6'b100011;
	  #10;
	  pressureData=6'b100100;
	  #10;
	  pressureData=6'b100101;
	  #10;
	  pressureData=6'b100110;
	  #10;
	  pressureData=6'b100111;
	  #10;
	  pressureData=6'b101000;
	  #10;
	  pressureData=6'b101001;
	  #10;
	  pressureData=6'b101010;
	  #10;
	  pressureData=6'b101011;
	  #10;
	  pressureData=6'b101100;
	  #10;
	  pressureData=6'b101101;
	  #10;
	  pressureData=6'b101110;
	  #10;
	  pressureData=6'b101111;
	  #10;
	  pressureData=6'b110000;
	  #10;
	  pressureData=6'b110001;
	  #10;
	  pressureData=6'b110010;
	  #10;
	  pressureData=6'b110011;
	  #10;
	  pressureData=6'b110100;
	  #10;
	  pressureData=6'b110101;
	  #10;
	  pressureData=6'b110110;
	  #10;
	  pressureData=6'b110111;
	  #10;
	  pressureData=6'b111000;
	  #10;
	  pressureData=6'b111001;
	  #10;
	  pressureData=6'b111010;
	  #10;
	  pressureData=6'b111011;
	  #10;
	  pressureData=6'b111100;
	  #10;
	  pressureData=6'b111101;
	  #10;
	  pressureData=6'b111110;
	  #10;
	  pressureData=6'b111111;
	  #10
	  bloodType <= 3'b000;
		# 5 ;
	   bloodPH <= 4'b0000;
		# 5 ;
		bloodPH <= 4'b0001;
		# 5 ;
		bloodPH <= 4'b0010;
		# 5 ;
		bloodPH <= 4'b0011;
		# 5 ;
		bloodPH <= 4'b0100;
		# 5 ;
		bloodPH <= 4'b0101;
		# 5 ;
		bloodPH <= 4'b0110;
		# 5 ;
		bloodPH <= 4'b0111;
		# 5 ;
		bloodPH <= 4'b1000;
		# 5 ;
		bloodPH <= 4'b1001;
		# 5 ;
		bloodPH <= 4'b1010;
		# 5 ;
		bloodPH <= 4'b1011;
		# 5 ;
		bloodPH <= 4'b1100;
		# 5 ;
		bloodPH <= 4'b1101;
		# 5 ;
		bloodPH <= 4'b1110;
		# 5 ;
		bloodPH <= 4'b1111;
		#10;
		bloodType <= 3'b001;
		# 5 ;
		bloodPH <= 4'b0000;
		# 5 ;
		bloodPH <= 4'b0001;
		# 5 ;
		bloodPH <= 4'b0010;
		# 5 ;
		bloodPH <= 4'b0011;
		# 5 ;
		bloodPH <= 4'b0100;
		# 5 ;
		bloodPH <= 4'b0101;
		# 5 ;
		bloodPH <= 4'b0110;
		# 5 ;
		bloodPH <= 4'b0111;
		# 5 ;
		bloodPH <= 4'b1000;
		# 5 ;
		bloodPH <= 4'b1001;
		# 5 ;
		bloodPH <= 4'b1010;
		# 5 ;
		bloodPH <= 4'b1011;
		# 5 ;
		bloodPH <= 4'b1100;
		# 5 ;
		bloodPH <= 4'b1101;
		# 5 ;
		bloodPH <= 4'b1110;
		# 5 ;
		bloodPH <= 4'b1111;
		#10;
		bloodType <= 3'b010;
		# 5 ;
		bloodPH <= 4'b0000;
		# 5 ;
		bloodPH <= 4'b0001;
		# 5 ;
		bloodPH <= 4'b0010;
		# 5 ;
		bloodPH <= 4'b0011;
		# 5 ;
		bloodPH <= 4'b0100;
		# 5 ;
		bloodPH <= 4'b0101;
		# 5 ;
		bloodPH <= 4'b0110;
		# 5 ;
		bloodPH <= 4'b0111;
		# 5 ;
		bloodPH <= 4'b1000;
		# 5 ;
		bloodPH <= 4'b1001;
		# 5 ;
		bloodPH <= 4'b1010;
		# 5 ;
		bloodPH <= 4'b1011;
		# 5 ;
		bloodPH <= 4'b1100;
		# 5 ;
		bloodPH <= 4'b1101;
		# 5 ;
		bloodPH <= 4'b1110;
		# 5 ;
		bloodPH <= 4'b1111;
		#10;
		bloodType <= 3'b011;
		# 5 ;
		bloodPH <= 4'b0000;
		# 5 ;
		bloodPH <= 4'b0001;
		# 5 ;
		bloodPH <= 4'b0010;
		# 5 ;
		bloodPH <= 4'b0011;
		# 5 ;
		bloodPH <= 4'b0100;
		# 5 ;
		bloodPH <= 4'b0101;
		# 5 ;
		bloodPH <= 4'b0110;
		# 5 ;
		bloodPH <= 4'b0111;
		# 5 ;
		bloodPH <= 4'b1000;
		# 5 ;
		bloodPH <= 4'b1001;
		# 5 ;
		bloodPH <= 4'b1010;
		# 5 ;
		bloodPH <= 4'b1011;
		# 5 ;
		bloodPH <= 4'b1100;
		# 5 ;
		bloodPH <= 4'b1101;
		# 5 ;
		bloodPH <= 4'b1110;
		# 5 ;
		bloodPH <= 4'b1111;
		#10;
		bloodType <= 3'b100;
		# 5 ;
		bloodPH <= 4'b0000;
		# 5 ;
		bloodPH <= 4'b0001;
		# 5 ;
		bloodPH <= 4'b0010;
		# 5 ;
		bloodPH <= 4'b0011;
		# 5 ;
		bloodPH <= 4'b0100;
		# 5 ;
		bloodPH <= 4'b0101;
		# 5 ;
		bloodPH <= 4'b0110;
		# 5 ;
		bloodPH <= 4'b0111;
		# 5 ;
		bloodPH <= 4'b1000;
		# 5 ;
		bloodPH <= 4'b1001;
		# 5 ;
		bloodPH <= 4'b1010;
		# 5 ;
		bloodPH <= 4'b1011;
		# 5 ;
		bloodPH <= 4'b1100;
		# 5 ;
		bloodPH <= 4'b1101;
		# 5 ;
		bloodPH <= 4'b1110;
		# 5 ;
		bloodPH <= 4'b1111;
		#10;
		bloodType <= 3'b101;
		# 5 ;
		bloodPH <= 4'b0000;
		# 5 ;
		bloodPH <= 4'b0001;
		# 5 ;
		bloodPH <= 4'b0010;
		# 5 ;
		bloodPH <= 4'b0011;
		# 5 ;
		bloodPH <= 4'b0100;
		# 5 ;
		bloodPH <= 4'b0101;
		# 5 ;
		bloodPH <= 4'b0110;
		# 5 ;
		bloodPH <= 4'b0111;
		# 5 ;
		bloodPH <= 4'b1000;
		# 5 ;
		bloodPH <= 4'b1001;
		# 5 ;
		bloodPH <= 4'b1010;
		# 5 ;
		bloodPH <= 4'b1011;
		# 5 ;
		bloodPH <= 4'b1100;
		# 5 ;
		bloodPH <= 4'b1101;
		# 5 ;
		bloodPH <= 4'b1110;
		# 5 ;
		bloodPH <= 4'b1111;
		#10;
		bloodType <= 3'b110;
		# 5 ;
		bloodPH <= 4'b0000;
		# 5 ;
		bloodPH <= 4'b0001;
		# 5 ;
		bloodPH <= 4'b0010;
		# 5 ;
		bloodPH <= 4'b0011;
		# 5 ;
		bloodPH <= 4'b0100;
		# 5 ;
		bloodPH <= 4'b0101;
		# 5 ;
		bloodPH <= 4'b0110;
		# 5 ;
		bloodPH <= 4'b0111;
		# 5 ;
		bloodPH <= 4'b1000;
		# 5 ;
		bloodPH <= 4'b1001;
		# 5 ;
		bloodPH <= 4'b1010;
		# 5 ;
		bloodPH <= 4'b1011;
		# 5 ;
		bloodPH <= 4'b1100;
		# 5 ;
		bloodPH <= 4'b1101;
		# 5 ;
		bloodPH <= 4'b1110;
		# 5 ;
		bloodPH <= 4'b1111;
		#10;
		bloodType <= 3'b111;
		# 5 ;
	   bloodPH <= 4'b0000;
		# 5 ;
		bloodPH <= 4'b0001;
		# 5 ;
		bloodPH <= 4'b0010;
		# 5 ;
		bloodPH <= 4'b0011;
		# 5 ;
		bloodPH <= 4'b0100;
		# 5 ;
		bloodPH <= 4'b0101;
		# 5 ;
		bloodPH <= 4'b0110;
		# 5 ;
		bloodPH <= 4'b0111;
		# 5 ;
		bloodPH <= 4'b1000;
		# 5 ;
		bloodPH <= 4'b1001;
		# 5 ;
		bloodPH <= 4'b1010;
		# 5 ;
		bloodPH <= 4'b1011;
		# 5 ;
		bloodPH <= 4'b1100;
		# 5 ;
		bloodPH <= 4'b1101;
		# 5 ;
		bloodPH <= 4'b1110;
		# 5 ;
		bloodPH <= 4'b1111;
		#10;
		fdFactoryValue = 8'b00010000;
		fdSensorValue= 8'b00000000;
		#5;
		fdSensorValue= 8'b00000001;
		#5;
		fdSensorValue= 8'b00000010;
		#5;
		fdSensorValue= 8'b00000011;
		#5;
		fdSensorValue= 8'b00000100;
		#5;
		fdSensorValue= 8'b00000101;
		#5;
		fdSensorValue= 8'b00000110;
		#5;
		fdSensorValue= 8'b00000111;
		#5;
		fdSensorValue= 8'b00001000;
		#5;
		fdSensorValue= 8'b00001001;
		#5;
		fdSensorValue= 8'b00001010;
		#5;
		fdSensorValue= 8'b00001011;
		#5;
		fdSensorValue= 8'b00001100;
		#5;
		fdSensorValue= 8'b00001101;
		#5;
		fdSensorValue= 8'b00001110;
		#5;
		fdSensorValue= 8'b00001111;
		#5;
		fdSensorValue= 8'b00010000;
		#5;
		fdSensorValue= 8'b00010001;
		#5;
		fdSensorValue= 8'b00010010;
		#5;
		fdSensorValue= 8'b00010011;
		#5;
		fdSensorValue= 8'b00010100;
		#5;
		fdSensorValue= 8'b00010101;
		#5;
		fdSensorValue= 8'b00010110;
		#5;
		fdSensorValue= 8'b00010111;
		#5;
		fdSensorValue= 8'b00011000;
		#5;
		fdSensorValue= 8'b00011001;
		#5;
		fdSensorValue= 8'b00011010;
		#5;
		fdSensorValue= 8'b00011011;
		#5;
		fdSensorValue= 8'b00011100;
		#5;
		fdSensorValue= 8'b00011101;
		#5;
		fdSensorValue= 8'b00011110;
		#5;
		fdSensorValue= 8'b00011111;
		#5;
		fdSensorValue= 8'b00100000;
		#5;
		fdSensorValue= 8'b00100001;
		#5;
		fdSensorValue= 8'b00100010;
		#5;
		fdSensorValue= 8'b00100011;
		#5;
		fdSensorValue= 8'b00100100;
		#5;
		fdSensorValue= 8'b00100101;
		#5;
		fdSensorValue= 8'b00100110;
		#5;
		fdSensorValue= 8'b00100111;
		#5;
		fdSensorValue= 8'b00101000;
		#5;
		fdSensorValue= 8'b00101001;
		#5;
		fdSensorValue= 8'b00101010;
		#5;
		fdSensorValue= 8'b00101011;
		#5;
		fdSensorValue= 8'b00101100;
		#5;
		fdSensorValue= 8'b00101101;
		#5;
		fdSensorValue= 8'b00101110;
		#5;
		fdSensorValue= 8'b00101111;
		#5;
		fdSensorValue= 8'b00110000;
		#5;
		fdSensorValue= 8'b00110001;
		#5;
		fdSensorValue= 8'b00110010;
		#5;
		fdSensorValue= 8'b00110011;
		#5;
		fdSensorValue= 8'b00110100;
		#5;
		fdSensorValue= 8'b00110101;
		#5;
		fdSensorValue= 8'b00110110;
		#5;
		fdSensorValue= 8'b00110111;
		#5;
		fdSensorValue= 8'b00111000;
		#5;
		fdSensorValue= 8'b00111001;
		#5;
		fdSensorValue= 8'b00111010;
		#5;
		fdSensorValue= 8'b00111011;
		#5;
		fdSensorValue= 8'b00111100;
		#5;
		fdSensorValue= 8'b00111101;
		#5;
		fdSensorValue= 8'b00111110;
		#5;
		fdSensorValue= 8'b00111111;
		#5;
		fdSensorValue= 8'b01000000;
		#5;
		fdSensorValue= 8'b01000001;
		#5;
		fdSensorValue= 8'b01000010;
		#5;
		fdSensorValue= 8'b01000011;
		#5;
		fdSensorValue= 8'b01000100;
		#5;
		fdSensorValue= 8'b01000101;
		#5;
		fdSensorValue= 8'b01000110;
		#5;
		fdSensorValue= 8'b01000111;
		#5;
		fdSensorValue= 8'b01001000;
		#5;
		fdSensorValue= 8'b01001001;
		#5;
		fdSensorValue= 8'b01001010;
		#5;
		fdSensorValue= 8'b01001011;
		#5;
		fdSensorValue= 8'b01001100;
		#5;
		fdSensorValue= 8'b01001101;
		#5;
		fdSensorValue= 8'b01001110;
		#5;
		fdSensorValue= 8'b01001111;
		#5;
		fdSensorValue= 8'b01010000;
		#5;
		fdSensorValue= 8'b01010001;
		#5;
		fdSensorValue= 8'b01010010;
		#5;
		fdSensorValue= 8'b01010011;
		#5;
		fdSensorValue= 8'b01010100;
		#5;
		fdSensorValue= 8'b01010101;
		#5;
		fdSensorValue= 8'b01010110;
		#5;
		fdSensorValue= 8'b01010111;
		#5;
		fdSensorValue= 8'b01011000;
		#5;
		fdSensorValue= 8'b01011001;
		#5;
		fdSensorValue= 8'b01011010;
		#5;
		fdSensorValue= 8'b01011011;
		#5;
		fdSensorValue= 8'b01011100;
		#5;
		fdSensorValue= 8'b01011101;
		#5;
		fdSensorValue= 8'b01011110;
		#5;
		fdSensorValue= 8'b01011111;
		#5;
		fdSensorValue= 8'b01100000;
		#5;
		fdSensorValue= 8'b01100001;
		#5;
		fdSensorValue= 8'b01100010;
		#5;
		fdSensorValue= 8'b01100011;
		#5;
		fdSensorValue= 8'b01100100;
		#5;
		fdSensorValue= 8'b01100101;
		#5;
		fdSensorValue= 8'b01100110;
		#5;
		fdSensorValue= 8'b01100111;
		#5;
		fdSensorValue= 8'b01101000;
		#5;
		fdSensorValue= 8'b01101001;
		#5;
		fdSensorValue= 8'b01101010;
		#5;
		fdSensorValue= 8'b01101011;
		#5;
		fdSensorValue= 8'b01101100;
		#5;
		fdSensorValue= 8'b01101101;
		#5;
		fdSensorValue= 8'b01101110;
		#5;
		fdSensorValue= 8'b01101111;
		#5;
		fdSensorValue= 8'b01110000;
		#5;
		fdSensorValue= 8'b01110001;
		#5;
		fdSensorValue= 8'b01110010;
		#5;
		fdSensorValue= 8'b01110011;
		#5;
		fdSensorValue= 8'b01110100;
		#5;
		fdSensorValue= 8'b01110101;
		#5;
		fdSensorValue= 8'b01110110;
		#5;
		fdSensorValue= 8'b01110111;
		#5;
		fdSensorValue= 8'b01111000;
		#5;
		fdSensorValue= 8'b01111001;
		#5;
		fdSensorValue= 8'b01111010;
		#5;
		fdSensorValue= 8'b01111011;
		#5;
		fdSensorValue= 8'b01111100;
		#5;
		fdSensorValue= 8'b01111101;
		#5;
		fdSensorValue= 8'b01111110;
		#5;
		fdSensorValue= 8'b01111111;
		#5;
		fdSensorValue= 8'b10000000;
		#5;
		fdSensorValue= 8'b10000001;
		#5;
		fdSensorValue= 8'b10000010;
		#5;
		fdSensorValue= 8'b10000011;
		#5;
		fdSensorValue= 8'b10000100;
		#5;
		fdSensorValue= 8'b10000101;
		#5;
		fdSensorValue= 8'b10000110;
		#5;
		fdSensorValue= 8'b10000111;
		#5;
		fdSensorValue= 8'b10001000;
		#5;
		fdSensorValue= 8'b10001001;
		#5;
		fdSensorValue= 8'b10001010;
		#5;
		fdSensorValue= 8'b10001011;
		#5;
		fdSensorValue= 8'b10001100;
		#5;
		fdSensorValue= 8'b10001101;
		#5;
		fdSensorValue= 8'b10001110;
		#5;
		fdSensorValue= 8'b10001111;
		#5;
		fdSensorValue= 8'b10010000;
		#5;
		fdSensorValue= 8'b10010001;
		#5;
		fdSensorValue= 8'b10010010;
		#5;
		fdSensorValue= 8'b10010011;
		#5;
		fdSensorValue= 8'b10010100;
		#5;
		fdSensorValue= 8'b10010101;
		#5;
		fdSensorValue= 8'b10010110;
		#5;
		fdSensorValue= 8'b10010111;
		#5;
		fdSensorValue= 8'b10011000;
		#5;
		fdSensorValue= 8'b10011001;
		#5;
		fdSensorValue= 8'b10011010;
		#5;
		fdSensorValue= 8'b10011011;
		#5;
		fdSensorValue= 8'b10011100;
		#5;
		fdSensorValue= 8'b10011101;
		#5;
		fdSensorValue= 8'b10011110;
		#5;
		fdSensorValue= 8'b10011111;
		#5;
		fdSensorValue= 8'b10100000;
		#5;
		fdSensorValue= 8'b10100001;
		#5;
		fdSensorValue= 8'b10100010;
		#5;
		fdSensorValue= 8'b10100011;
		#5;
		fdSensorValue= 8'b10100100;
		#5;
		fdSensorValue= 8'b10100101;
		#5;
		fdSensorValue= 8'b10100110;
		#5;
		fdSensorValue= 8'b10100111;
		#5;
		fdSensorValue= 8'b10101000;
		#5;
		fdSensorValue= 8'b10101001;
		#5;
		fdSensorValue= 8'b10101010;
		#5;
		fdSensorValue= 8'b10101011;
		#5;
		fdSensorValue= 8'b10101100;
		#5;
		fdSensorValue= 8'b10101101;
		#5;
		fdSensorValue= 8'b10101110;
		#5;
		fdSensorValue= 8'b10101111;
		#5;
		fdSensorValue= 8'b10110000;
		#5;
		fdSensorValue= 8'b10110001;
		#5;
		fdSensorValue= 8'b10110010;
		#5;
		fdSensorValue= 8'b10110011;
		#5;
		fdSensorValue= 8'b10110100;
		#5;
		fdSensorValue= 8'b10110101;
		#5;
		fdSensorValue= 8'b10110110;
		#5;
		fdSensorValue= 8'b10110111;
		#5;
		fdSensorValue= 8'b10111000;
		#5;
		fdSensorValue= 8'b10111001;
		#5;
		fdSensorValue= 8'b10111010;
		#5;
		fdSensorValue= 8'b10111011;
		#5;
		fdSensorValue= 8'b10111100;
		#5;
		fdSensorValue= 8'b10111101;
		#5;
		fdSensorValue= 8'b10111110;
		#5;
		fdSensorValue= 8'b10111111;
		#5;
		fdSensorValue= 8'b11000000;
		#5;
		fdSensorValue= 8'b11000001;
		#5;
		fdSensorValue= 8'b11000010;
		#5;
		fdSensorValue= 8'b11000011;
		#5;
		fdSensorValue= 8'b11000100;
		#5;
		fdSensorValue= 8'b11000101;
		#5;
		fdSensorValue= 8'b11000110;
		#5;
		fdSensorValue= 8'b11000111;
		#5;
		fdSensorValue= 8'b11001000;
		#5;
		fdSensorValue= 8'b11001001;
		#5;
		fdSensorValue= 8'b11001010;
		#5;
		fdSensorValue= 8'b11001011;
		#5;
		fdSensorValue= 8'b11001100;
		#5;
		fdSensorValue= 8'b11001101;
		#5;
		fdSensorValue= 8'b11001110;
		#5;
		fdSensorValue= 8'b11001111;
		#5;
		fdSensorValue= 8'b11010000;
		#5;
		fdSensorValue= 8'b11010001;
		#5;
		fdSensorValue= 8'b11010010;
		#5;
		fdSensorValue= 8'b11010011;
		#5;
		fdSensorValue= 8'b11010100;
		#5;
		fdSensorValue= 8'b11010101;
		#5;
		fdSensorValue= 8'b11010110;
		#5;
		fdSensorValue= 8'b11010111;
		#5;
		fdSensorValue= 8'b11011000;
		#5;
		fdSensorValue= 8'b11011001;
		#5;
		fdSensorValue= 8'b11011010;
		#5;
		fdSensorValue= 8'b11011011;
		#5;
		fdSensorValue= 8'b11011100;
		#5;
		fdSensorValue= 8'b11011101;
		#5;
		fdSensorValue= 8'b11011110;
		#5;
		fdSensorValue= 8'b11011111;
		#5;
		fdSensorValue= 8'b11100000;
		#5;
		fdSensorValue= 8'b11100001;
		#5;
		fdSensorValue= 8'b11100010;
		#5;
		fdSensorValue= 8'b11100011;
		#5;
		fdSensorValue= 8'b11100100;
		#5;
		fdSensorValue= 8'b11100101;
		#5;
		fdSensorValue= 8'b11100110;
		#5;
		fdSensorValue= 8'b11100111;
		#5;
		fdSensorValue= 8'b11101000;
		#5;
		fdSensorValue= 8'b11101001;
		#5;
		fdSensorValue= 8'b11101010;
		#5;
		fdSensorValue= 8'b11101011;
		#5;
		fdSensorValue= 8'b11101100;
		#5;
		fdSensorValue= 8'b11101101;
		#5;
		fdSensorValue= 8'b11101110;
		#5;
		fdSensorValue= 8'b11101111;
		#5;
		fdSensorValue= 8'b11110000;
		#5;
		fdSensorValue= 8'b11110001;
		#5;
		fdSensorValue= 8'b11110010;
		#5;
		fdSensorValue= 8'b11110011;
		#5;
		fdSensorValue= 8'b11110100;
		#5;
		fdSensorValue= 8'b11110101;
		#5;
		fdSensorValue= 8'b11110110;
		#5;
		fdSensorValue= 8'b11110111;
		#5;
		fdSensorValue= 8'b11111000;
		#5;
		fdSensorValue= 8'b11111001;
		#5;
		fdSensorValue= 8'b11111010;
		#5;
		fdSensorValue= 8'b11111011;
		#5;
		fdSensorValue= 8'b11111100;
		#5;
		fdSensorValue= 8'b11111101;
		#5;
		fdSensorValue= 8'b11111110;
		#5;
		fdSensorValue= 8'b11111111;
		#5;
		factotyBaseTemp <= 5'b00001;
      factotyTempCoef <= 4'b1000;
		tempSensorValue <= 4'b0000;
		# 10 ;
		tempSensorValue <= 4'b0001;
		# 10;
	   tempSensorValue <= 4'b0010;
		# 10;
		tempSensorValue <=4'b0011;
		# 10 ;
		tempSensorValue <=4'b0100;
		# 10 ;
	   tempSensorValue <= 4'b0101;
		# 10;
		tempSensorValue <=4'b0110;
		# 10 ;
	   tempSensorValue <= 4'b0111;
		# 10;
		tempSensorValue <=4'b1000;
		# 10 ;
	   tempSensorValue <= 4'b1001;
		# 10;
		tempSensorValue <=4'b1010;
		# 10 ;
	   tempSensorValue <= 4'b1011;
		# 10;
		tempSensorValue <=4'b1100;		
	   # 10 ;
		tempSensorValue <=4'b1101;
		# 10 ;
		tempSensorValue <=4'b1110;
		# 10 ;
		tempSensorValue <=4'b1111;
		# 10 ;
		bloodSensor = 8'b00000000;
		#5;
		bloodSensor = 8'b00000001;
		#5;
		bloodSensor = 8'b00000010;
		#5;
		bloodSensor = 8'b00000011;
		#5;
		bloodSensor = 8'b00000100;
		#5;
		bloodSensor = 8'b00000101;
		#5;
		bloodSensor = 8'b00000110;
		#5;
		bloodSensor = 8'b00000111;
		#5;
		bloodSensor = 8'b00001000;
		#5;
		bloodSensor = 8'b00001001;
		#5;
		bloodSensor = 8'b00001010;
		#5;
		bloodSensor = 8'b00001011;
		#5;
		bloodSensor = 8'b00001100;
		#5;
		bloodSensor = 8'b00001101;
		#5;
		bloodSensor = 8'b00001110;
		#5;
		bloodSensor = 8'b00001111;
		#5;
		bloodSensor = 8'b00010000;
		#5;
		bloodSensor = 8'b00010001;
		#5;
		bloodSensor = 8'b00010010;
		#5;
		bloodSensor = 8'b00010011;
		#5;
		bloodSensor = 8'b00010100;
		#5;
		bloodSensor = 8'b00010101;
		#5;
		bloodSensor = 8'b00010110;
		#5;
		bloodSensor = 8'b00010111;
		#5;
		bloodSensor = 8'b00011000;
		#5;
		bloodSensor = 8'b00011001;
		#5;
		bloodSensor = 8'b00011010;
		#5;
		bloodSensor = 8'b00011011;
		#5;
		bloodSensor = 8'b00011100;
		#5;
		bloodSensor = 8'b00011101;
		#5;
		bloodSensor = 8'b00011110;
		#5;
		bloodSensor = 8'b00011111;
		#5;
		bloodSensor = 8'b00100000;
		#5;
		bloodSensor = 8'b00100001;
		#5;
		bloodSensor = 8'b00100010;
		#5;
		bloodSensor = 8'b00100011;
		#5;
		bloodSensor = 8'b00100100;
		#5;
		bloodSensor = 8'b00100101;
		#5;
		bloodSensor = 8'b00100110;
		#5;
		bloodSensor = 8'b00100111;
		#5;
		bloodSensor = 8'b00101000;
		#5;
		bloodSensor = 8'b00101001;
		#5;
		bloodSensor = 8'b00101010;
		#5;
		bloodSensor = 8'b00101011;
		#5;
		bloodSensor = 8'b00101100;
		#5;
		bloodSensor = 8'b00101101;
		#5;
		bloodSensor = 8'b00101110;
		#5;
		bloodSensor = 8'b00101111;
		#5;
		bloodSensor = 8'b00110000;
		#5;
		bloodSensor = 8'b00110001;
		#5;
		bloodSensor = 8'b00110010;
		#5;
		bloodSensor = 8'b00110011;
		#5;
		bloodSensor = 8'b00110100;
		#5;
		bloodSensor = 8'b00110101;
		#5;
		bloodSensor = 8'b00110110;
		#5;
		bloodSensor = 8'b00110111;
		#5;
		bloodSensor = 8'b00111000;
		#5;
		bloodSensor = 8'b00111001;
		#5;
		bloodSensor = 8'b00111010;
		#5;
		bloodSensor = 8'b00111011;
		#5;
		bloodSensor = 8'b00111100;
		#5;
		bloodSensor = 8'b00111101;
		#5;
		bloodSensor = 8'b00111110;
		#5;
		bloodSensor = 8'b00111111;
		#5;
		bloodSensor = 8'b01000000;
		#5;
		bloodSensor = 8'b01000001;
		#5;
		bloodSensor = 8'b01000010;
		#5;
		bloodSensor = 8'b01000011;
		#5;
		bloodSensor = 8'b01000100;
		#5;
		bloodSensor = 8'b01000101;
		#5;
		bloodSensor = 8'b01000110;
		#5;
		bloodSensor = 8'b01000111;
		#5;
		bloodSensor = 8'b01001000;
		#5;
		bloodSensor = 8'b01001001;
		#5;
		bloodSensor = 8'b01001010;
		#5;
		bloodSensor = 8'b01001011;
		#5;
		bloodSensor = 8'b01001100;
		#5;
		bloodSensor = 8'b01001101;
		#5;
		bloodSensor = 8'b01001110;
		#5;
		bloodSensor = 8'b01001111;
		#5;
		bloodSensor = 8'b01010000;
		#5;
		bloodSensor = 8'b01010001;
		#5;
		bloodSensor = 8'b01010010;
		#5;
		bloodSensor = 8'b01010011;
		#5;
		bloodSensor = 8'b01010100;
		#5;
		bloodSensor = 8'b01010101;
		#5;
		bloodSensor = 8'b01010110;
		#5;
		bloodSensor = 8'b01010111;
		#5;
		bloodSensor = 8'b01011000;
		#5;
		bloodSensor = 8'b01011001;
		#5;
		bloodSensor = 8'b01011010;
		#5;
		bloodSensor = 8'b01011011;
		#5;
		bloodSensor = 8'b01011100;
		#5;
		bloodSensor = 8'b01011101;
		#5;
		bloodSensor = 8'b01011110;
		#5;
		bloodSensor = 8'b01011111;
		#5;
		bloodSensor = 8'b01100000;
		#5;
		bloodSensor = 8'b01100001;
		#5;
		bloodSensor = 8'b01100010;
		#5;
		bloodSensor = 8'b01100011;
		#5;
		bloodSensor = 8'b01100100;
		#5;
		bloodSensor = 8'b01100101;
		#5;
		bloodSensor = 8'b01100110;
		#5;
		bloodSensor = 8'b01100111;
		#5;
		bloodSensor = 8'b01101000;
		#5;
		bloodSensor = 8'b01101001;
		#5;
		bloodSensor = 8'b01101010;
		#5;
		bloodSensor = 8'b01101011;
		#5;
		bloodSensor = 8'b01101100;
		#5;
		bloodSensor = 8'b01101101;
		#5;
		bloodSensor = 8'b01101110;
		#5;
		bloodSensor = 8'b01101111;
		#5;
		bloodSensor = 8'b01110000;
		#5;
		bloodSensor = 8'b01110001;
		#5;
		bloodSensor = 8'b01110010;
		#5;
		bloodSensor = 8'b01110011;
		#5;
		bloodSensor = 8'b01110100;
		#5;
		bloodSensor = 8'b01110101;
		#5;
		bloodSensor = 8'b01110110;
		#5;
		bloodSensor = 8'b01110111;
		#5;
		bloodSensor = 8'b01111000;
		#5;
		bloodSensor = 8'b01111001;
		#5;
		bloodSensor = 8'b01111010;
		#5;
		bloodSensor = 8'b01111011;
		#5;
		bloodSensor = 8'b01111100;
		#5;
		bloodSensor = 8'b01111101;
		#5;
		bloodSensor = 8'b01111110;
		#5;
		bloodSensor = 8'b01111111;
		#5;
		bloodSensor = 8'b10000000;
		#5;
		bloodSensor = 8'b10000001;
		#5;
		bloodSensor = 8'b10000010;
		#5;
		bloodSensor = 8'b10000011;
		#5;
		bloodSensor = 8'b10000100;
		#5;
		bloodSensor = 8'b10000101;
		#5;
		bloodSensor = 8'b10000110;
		#5;
		bloodSensor = 8'b10000111;
		#5;
		bloodSensor = 8'b10001000;
		#5;
		bloodSensor = 8'b10001001;
		#5;
		bloodSensor = 8'b10001010;
		#5;
		bloodSensor = 8'b10001011;
		#5;
		bloodSensor = 8'b10001100;
		#5;
		bloodSensor = 8'b10001101;
		#5;
		bloodSensor = 8'b10001110;
		#5;
		bloodSensor = 8'b10001111;
		#5;
		bloodSensor = 8'b10010000;
		#5;
		bloodSensor = 8'b10010001;
		#5;
		bloodSensor = 8'b10010010;
		#5;
		bloodSensor = 8'b10010011;
		#5;
		bloodSensor = 8'b10010100;
		#5;
		bloodSensor = 8'b10010101;
		#5;
		bloodSensor = 8'b10010110;
		#5;
		bloodSensor = 8'b10010111;
		#5;
		bloodSensor = 8'b10011000;
		#5;
		bloodSensor = 8'b10011001;
		#5;
		bloodSensor = 8'b10011010;
		#5;
		bloodSensor = 8'b10011011;
		#5;
		bloodSensor = 8'b10011100;
		#5;
		bloodSensor = 8'b10011101;
		#5;
		bloodSensor = 8'b10011110;
		#5;
		bloodSensor = 8'b10011111;
		#5;
		bloodSensor = 8'b10100000;
		#5;
		bloodSensor = 8'b10100001;
		#5;
		bloodSensor = 8'b10100010;
		#5;
		bloodSensor = 8'b10100011;
		#5;
		bloodSensor = 8'b10100100;
		#5;
		bloodSensor = 8'b10100101;
		#5;
		bloodSensor = 8'b10100110;
		#5;
		bloodSensor = 8'b10100111;
		#5;
		bloodSensor = 8'b10101000;
		#5;
		bloodSensor = 8'b10101001;
		#5;
		bloodSensor = 8'b10101010;
		#5;
		bloodSensor = 8'b10101011;
		#5;
		bloodSensor = 8'b10101100;
		#5;
		bloodSensor = 8'b10101101;
		#5;
		bloodSensor = 8'b10101110;
		#5;
		bloodSensor = 8'b10101111;
		#5;
		bloodSensor = 8'b10110000;
		#5;
		bloodSensor = 8'b10110001;
		#5;
		bloodSensor = 8'b10110010;
		#5;
		bloodSensor = 8'b10110011;
		#5;
		bloodSensor = 8'b10110100;
		#5;
		bloodSensor = 8'b10110101;
		#5;
		bloodSensor = 8'b10110110;
		#5;
		bloodSensor = 8'b10110111;
		#5;
		bloodSensor = 8'b10111000;
		#5;
		bloodSensor = 8'b10111001;
		#5;
		bloodSensor = 8'b10111010;
		#5;
		bloodSensor = 8'b10111011;
		#5;
		bloodSensor = 8'b10111100;
		#5;
		bloodSensor = 8'b10111101;
		#5;
		bloodSensor = 8'b10111110;
		#5;
		bloodSensor = 8'b10111111;
		#5;
		bloodSensor = 8'b11000000;
		#5;
		bloodSensor = 8'b11000001;
		#5;
		bloodSensor = 8'b11000010;
		#5;
		bloodSensor = 8'b11000011;
		#5;
		bloodSensor = 8'b11000100;
		#5;
		bloodSensor = 8'b11000101;
		#5;
		bloodSensor = 8'b11000110;
		#5;
		bloodSensor = 8'b11000111;
		#5;
		bloodSensor = 8'b11001000;
		#5;
		bloodSensor = 8'b11001001;
		#5;
		bloodSensor = 8'b11001010;
		#5;
		bloodSensor = 8'b11001011;
		#5;
		bloodSensor = 8'b11001100;
		#5;
		bloodSensor = 8'b11001101;
		#5;
		bloodSensor = 8'b11001110;
		#5;
		bloodSensor = 8'b11001111;
		#5;
		bloodSensor = 8'b11010000;
		#5;
		bloodSensor = 8'b11010001;
		#5;
		bloodSensor = 8'b11010010;
		#5;
		bloodSensor = 8'b11010011;
		#5;
		bloodSensor = 8'b11010100;
		#5;
		bloodSensor = 8'b11010101;
		#5;
		bloodSensor = 8'b11010110;
		#5;
		bloodSensor = 8'b11010111;
		#5;
		bloodSensor = 8'b11011000;
		#5;
		bloodSensor = 8'b11011001;
		#5;
		bloodSensor = 8'b11011010;
		#5;
		bloodSensor = 8'b11011011;
		#5;
		bloodSensor = 8'b11011100;
		#5;
		bloodSensor = 8'b11011101;
		#5;
		bloodSensor = 8'b11011110;
		#5;
		bloodSensor = 8'b11011111;
		#5;
		bloodSensor = 8'b11100000;
		#5;
		bloodSensor = 8'b11100001;
		#5;
		bloodSensor = 8'b11100010;
		#5;
		bloodSensor = 8'b11100011;
		#5;
		bloodSensor = 8'b11100100;
		#5;
		bloodSensor = 8'b11100101;
		#5;
		bloodSensor = 8'b11100110;
		#5;
		bloodSensor = 8'b11100111;
		#5;
		bloodSensor = 8'b11101000;
		#5;
		bloodSensor = 8'b11101001;
		#5;
		bloodSensor = 8'b11101010;
		#5;
		bloodSensor = 8'b11101011;
		#5;
		bloodSensor = 8'b11101100;
		#5;
		bloodSensor = 8'b11101101;
		#5;
		bloodSensor = 8'b11101110;
		#5;
		bloodSensor = 8'b11101111;
		#5;
		bloodSensor = 8'b11110000;
		#5;
		bloodSensor = 8'b11110001;
		#5;
		bloodSensor = 8'b11110010;
		#5;
		bloodSensor = 8'b11110011;
		#5;
		bloodSensor = 8'b11110100;
		#5;
		bloodSensor = 8'b11110101;
		#5;
		bloodSensor = 8'b11110110;
		#5;
		bloodSensor = 8'b11110111;
		#5;
		bloodSensor = 8'b11111000;
		#5;
		bloodSensor = 8'b11111001;
		#5;
		bloodSensor = 8'b11111010;
		#5;
		bloodSensor = 8'b11111011;
		#5;
		bloodSensor = 8'b11111100;
		#5;
		bloodSensor = 8'b11111101;
		#5;
		bloodSensor = 8'b11111110;
		#5;
		bloodSensor = 8'b11111111;
		#5;
		$finish;
	end

endmodule
